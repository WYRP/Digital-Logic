-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions
-- and other software and tools, and its AMPP partner logic
-- functions, and any output files from any of the foregoing
-- (including device programming or simulation files), and any
-- associated documentation or information are expressly subject
-- to the terms and conditions of the Altera Program License
-- Subscription Agreement, Altera MegaCore Function License
-- Agreement, or other applicable license agreement, including,
-- without limitation, that your use is for the sole purpose of
-- programming logic devices manufactured by Altera and sold by
-- Altera or its authorized distributors.  Please refer to the
-- applicable agreement for further details.

-- PROGRAM "Quartus II 64-Bit"
-- VERSION "Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED "Tue Feb 08 13:31:36 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY work;

ENTITY chenyi_xu_4bit_barrel IS
PORT
(
sel :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
X :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
Y :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
);
END chenyi_xu_4bit_barrel;

ARCHITECTURE bdf_type OF chenyi_xu_4bit_barrel IS

SIGNAL SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL SYNTHESIZED_WIRE_29 :  STD_LOGIC;


BEGIN



SYNTHESIZED_WIRE_2 <= SYNTHESIZED_WIRE_32 AND X(0);


SYNTHESIZED_WIRE_1 <= sel(1) AND X(2);


SYNTHESIZED_WIRE_34 <= SYNTHESIZED_WIRE_1 OR SYNTHESIZED_WIRE_2;


SYNTHESIZED_WIRE_36 <= SYNTHESIZED_WIRE_3 OR SYNTHESIZED_WIRE_4;


SYNTHESIZED_WIRE_37 <= SYNTHESIZED_WIRE_5 OR SYNTHESIZED_WIRE_6;


SYNTHESIZED_WIRE_35 <= SYNTHESIZED_WIRE_7 OR SYNTHESIZED_WIRE_8;


SYNTHESIZED_WIRE_23 <= SYNTHESIZED_WIRE_33 AND SYNTHESIZED_WIRE_34;


SYNTHESIZED_WIRE_22 <= sel(0) AND SYNTHESIZED_WIRE_35;


SYNTHESIZED_WIRE_25 <= SYNTHESIZED_WIRE_33 AND SYNTHESIZED_WIRE_36;


SYNTHESIZED_WIRE_24 <= sel(0) AND SYNTHESIZED_WIRE_34;


SYNTHESIZED_WIRE_4 <= SYNTHESIZED_WIRE_32 AND X(1);


SYNTHESIZED_WIRE_27 <= SYNTHESIZED_WIRE_33 AND SYNTHESIZED_WIRE_37;


SYNTHESIZED_WIRE_26 <= sel(0) AND SYNTHESIZED_WIRE_36;


SYNTHESIZED_WIRE_29 <= SYNTHESIZED_WIRE_33 AND SYNTHESIZED_WIRE_35;


SYNTHESIZED_WIRE_28 <= sel(0) AND SYNTHESIZED_WIRE_37;


Y(0) <= SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_23;


Y(1) <= SYNTHESIZED_WIRE_24 OR SYNTHESIZED_WIRE_25;


Y(2) <= SYNTHESIZED_WIRE_26 OR SYNTHESIZED_WIRE_27;


Y(3) <= SYNTHESIZED_WIRE_28 OR SYNTHESIZED_WIRE_29;


SYNTHESIZED_WIRE_3 <= sel(1) AND X(3);


SYNTHESIZED_WIRE_6 <= SYNTHESIZED_WIRE_32 AND X(0);


SYNTHESIZED_WIRE_5 <= sel(1) AND X(2);


SYNTHESIZED_WIRE_8 <= SYNTHESIZED_WIRE_32 AND X(1);


SYNTHESIZED_WIRE_7 <= sel(1) AND X(3);


SYNTHESIZED_WIRE_32 <= NOT(sel(1));



SYNTHESIZED_WIRE_33 <= NOT(sel(0));



END bdf_type;